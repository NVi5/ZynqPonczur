`timescale 1ns / 1ps
`include "bmp.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 04.05.2021 20:54:38
// Design Name:
// Module Name: behav_tb
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module behav_tb();
    integer vertices[] = {
        -19,19,-19,19,-19,-19,-19,-19,-19,19,-19,19,54,19,19,19,19,19,19,19,19,-19,-19,19,19,-19,19,-19,-19,-19,-199,19,-19,-19,19,-19,-19,-19,-19,-19,-123,19,-19,-19,19,19,19,19,-19,55,19,-19,19,19,-19,55,-19,19,95,-19,19,55,-19,-19,19,-19,19,55,-19,19,19,-19,-19,19,19,-19,55,-19,-19,19,-19,19,19,-19,19,55,19,19,19,19,19,95,-19,-19,95,19,19,95,19,-19,55,19,-19,95,-19,-19,55,-19,19,95,19,274,95,-19,19,95,-19,19,55,19,-19,95,19,-19,55,19,274,95,-19,313,55,-19,274,55,-19,19,55,-19,274,55,19,19,55,19,19,55,19,274,95,19,19,95,19,19,95,-19,274,55,-19,19,55,-19,313,55,-19,313,95,19,313,55,19,274,55,-19,313,55,19,274,55,19,274,55,19,313,95,19,274,95,19,313,95,19,274,151,19,274,95,19,274,151,19,313,151,-19,274,151,-19,313,95,-19,313,151,19,313,95,19,274,95,19,274,151,-19,274,95,-19,274,95,-19,313,151,-19,313,95,-19,-19,-123,19,19,-163,19,19,-123,19,19,-19,19,19,-123,-19,19,-19,-19,19,-19,-19,-19,-123,-19,-19,-19,-19,-19,-19,19,19,-123,19,19,-19,19,19,-163,19,-19,-163,-19,19,-163,-19,19,-123,-19,-19,-163,-19,-19,-123,-19,-19,-163,-19,-138,-123,-19,-19,-123,-19,19,-123,19,19,-163,-19,19,-123,-19,-138,-123,-19,-138,-163,19,-138,-123,19,-19,-163,19,-138,-163,-19,-19,-163,-19,-19,-123,-19,-138,-123,19,-19,-123,19,-19,-123,19,-138,-163,19,-19,-163,19,-199,-19,19,-199,-91,-19,-199,-19,-19,-19,-19,19,-199,-19,-19,-19,-19,-19,-19,19,-19,-199,19,19,-19,19,19,-19,19,19,-199,-19,19,-19,-19,19,-245,19,19,-245,-19,-19,-245,-19,19,-199,-19,-19,-245,19,-19,-199,19,-19,-199,19,-19,-245,19,19,-199,19,19,-199,19,19,-245,-19,19,-199,-19,19,-199,-91,19,-245,-91,-19,-199,-91,-19,-199,-19,-19,-245,-91,-19,-245,-19,-19,-245,-19,19,-199,-91,19,-199,-19,19,-245,-19,-19,-245,-91,19,-245,-19,19,54,19,-19,90,-19,-19,54,-19,-19,19,-19,-19,54,-19,19,19,-19,19,19,19,19,54,19,-19,19,19,-19,19,19,-19,54,-19,-19,19,-19,-19,90,19,-19,90,-19,19,90,-19,-19,54,-19,19,90,19,19,54,19,19,90,-19,19,90,-163,-19,90,-19,-19,54,19,19,90,19,-19,54,19,-19,90,-163,-19,54,-195,-19,54,-163,-19,54,-19,19,90,-163,19,90,-19,19,54,-19,-19,54,-163,19,54,-19,19,90,-19,-19,54,-163,-19,54,-19,-19,54,-195,-19,90,-195,19,54,-195,19,54,-163,-19,54,-195,19,54,-163,19,54,-163,19,90,-195,19,90,-163,19,90,-195,19,310,-163,19,90,-163,19,310,-163,19,310,-195,-19,310,-163,-19,90,-195,-19,310,-195,19,90,-195,19,90,-163,19,310,-163,-19,90,-163,-19,90,-163,-19,310,-195,-19,90,-195,-19,-19,19,-19,19,19,-19,19,-19,-19,19,-19,19,54,-19,19,54,19,19,19,19,19,-19,19,19,-19,-19,19,-19,-19,-19,-199,-19,-19,-199,19,-19,-19,-19,-19,-19,-123,-19,-19,-123,19,19,19,19,19,55,19,-19,55,19,-19,55,-19,-19,95,-19,19,95,-19,-19,19,-19,-19,55,-19,19,55,-19,-19,19,19,-19,55,19,-19,55,-19,19,19,-19,19,55,-19,19,55,19,19,95,-19,-19,95,-19,-19,95,19,-19,55,19,-19,95,19,-19,95,-19,19,95,19,274,95,19,274,95,-19,19,55,19,19,95,19,-19,95,19,274,95,-19,313,95,-19,313,55,-19,19,55,-19,274,55,-19,274,55,19,19,55,19,274,55,19,274,95,19,19,95,-19,274,95,-19,274,55,-19,313,55,-19,313,95,-19,313,95,19,274,55,-19,313,55,-19,313,55,19,274,55,19,313,55,19,313,95,19,313,95,19,313,151,19,274,151,19,274,151,19,313,151,19,313,151,-19,313,95,-19,313,151,-19,313,151,19,274,95,19,274,151,19,274,151,-19,274,95,-19,274,151,-19,313,151,-19,-19,-123,19,-19,-163,19,19,-163,19,19,-19,19,19,-123,19,19,-123,-19,19,-19,-19,19,-123,-19,-19,-123,-19,-19,-19,19,-19,-123,19,19,-123,19,19,-163,19,-19,-163,19,-19,-163,-19,19,-123,-19,19,-163,-19,-19,-163,-19,-19,-163,-19,-138,-163,-19,-138,-123,-19,19,-123,19,19,-163,19,19,-163,-19,-138,-123,-19,-138,-163,-19,-138,-163,19,-19,-163,19,-138,-163,19,-138,-163,-19,-19,-123,-19,-138,-123,-19,-138,-123,19,-19,-123,19,-138,-123,19,-138,-163,19,-199,-19,19,-199,-91,19,-199,-91,-19,-19,-19,19,-199,-19,19,-199,-19,-19,-19,19,-19,-199,19,-19,-199,19,19,-19,19,19,-199,19,19,-199,-19,19,-245,19,19,-245,19,-19,-245,-19,-19,-199,-19,-19,-245,-19,-19,-245,19,-19,-199,19,-19,-245,19,-19,-245,19,19,-199,19,19,-245,19,19,-245,-19,19,-199,-91,19,-245,-91,19,-245,-91,-19,-199,-19,-19,-199,-91,-19,-245,-91,-19,-245,-19,19,-245,-91,19,-199,-91,19,-245,-19,-19,-245,-91,-19,-245,-91,19,54,19,-19,90,19,-19,90,-19,-19,19,-19,-19,54,-19,-19,54,-19,19,19,19,19,54,19,19,54,19,-19,19,19,-19,54,19,-19,54,-19,-19,90,19,-19,90,19,19,90,-19,19,54,-19,19,90,-19,19,90,19,19,90,-19,19,90,-163,19,90,-163,-19,54,19,19,90,19,19,90,19,-19,90,-163,-19,90,-195,-19,54,-195,-19,54,-19,19,54,-163,19,90,-163,19,54,-19,-19,54,-163,-19,54,-163,19,90,-19,-19,90,-163,-19,54,-163,-19,54,-195,-19,90,-195,-19,90,-195,19,54,-163,-19,54,-195,-19,54,-195,19,54,-163,19,54,-195,19,90,-195,19,90,-195,19,310,-195,19,310,-163,19,310,-163,19,310,-195,19,310,-195,-19,90,-195,-19,310,-195,-19,310,-195,19,90,-163,19,310,-163,19,310,-163,-19,90,-163,-19,310,-163,-19,310,-195,-19
    };
    reg [7:0] framebuffer[800*600];

    rasterize_behav restarizer_i(vertices, framebuffer, $size(vertices));

    initial begin
        integer file;
        file = $fopen("picture.bmp", "wb");
        for (integer i=0;i<1078;i=i+1) begin
            $fwrite(file, "%c", bmp_header[i]);
        end
        for (integer y = 0; y < 600; y = y + 1) begin
            for (integer x = 0; x < 800; x = x + 1) begin
                $fwrite(file, "%c", framebuffer[y * 800 + x]);
            end
        end
        $fclose(file);
    end
endmodule

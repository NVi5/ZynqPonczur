`ifndef BMP_HEADER
`define BMP_HEADER

reg [7:0] bmp_header [0:1077] = {
    8'h42, 8'h4d, 8'h36, 8'h57, 8'h07, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h36, 8'h04,
    8'h00, 8'h00, 8'h28, 8'h00, 8'h00, 8'h00, 8'h20, 8'h03, 8'h00, 8'h00, 8'h58, 8'h02,
    8'h00, 8'h00, 8'h01, 8'h00, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53,
    8'h07, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h80, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h80, 8'h80, 8'h00, 8'h80, 8'h00,
    8'h00, 8'h00, 8'h80, 8'h00, 8'h80, 8'h00, 8'h80, 8'h80, 8'h00, 8'h00, 8'hc0, 8'hc0,
    8'hc0, 8'h00, 8'hc0, 8'hdc, 8'hc0, 8'h00, 8'hf0, 8'hca, 8'ha6, 8'h00, 8'h00, 8'h20,
    8'h40, 8'h00, 8'h00, 8'h20, 8'h60, 8'h00, 8'h00, 8'h20, 8'h80, 8'h00, 8'h00, 8'h20,
    8'ha0, 8'h00, 8'h00, 8'h20, 8'hc0, 8'h00, 8'h00, 8'h20, 8'he0, 8'h00, 8'h00, 8'h40,
    8'h00, 8'h00, 8'h00, 8'h40, 8'h20, 8'h00, 8'h00, 8'h40, 8'h40, 8'h00, 8'h00, 8'h40,
    8'h60, 8'h00, 8'h00, 8'h40, 8'h80, 8'h00, 8'h00, 8'h40, 8'ha0, 8'h00, 8'h00, 8'h40,
    8'hc0, 8'h00, 8'h00, 8'h40, 8'he0, 8'h00, 8'h00, 8'h60, 8'h00, 8'h00, 8'h00, 8'h60,
    8'h20, 8'h00, 8'h00, 8'h60, 8'h40, 8'h00, 8'h00, 8'h60, 8'h60, 8'h00, 8'h00, 8'h60,
    8'h80, 8'h00, 8'h00, 8'h60, 8'ha0, 8'h00, 8'h00, 8'h60, 8'hc0, 8'h00, 8'h00, 8'h60,
    8'he0, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h80, 8'h20, 8'h00, 8'h00, 8'h80,
    8'h40, 8'h00, 8'h00, 8'h80, 8'h60, 8'h00, 8'h00, 8'h80, 8'h80, 8'h00, 8'h00, 8'h80,
    8'ha0, 8'h00, 8'h00, 8'h80, 8'hc0, 8'h00, 8'h00, 8'h80, 8'he0, 8'h00, 8'h00, 8'ha0,
    8'h00, 8'h00, 8'h00, 8'ha0, 8'h20, 8'h00, 8'h00, 8'ha0, 8'h40, 8'h00, 8'h00, 8'ha0,
    8'h60, 8'h00, 8'h00, 8'ha0, 8'h80, 8'h00, 8'h00, 8'ha0, 8'ha0, 8'h00, 8'h00, 8'ha0,
    8'hc0, 8'h00, 8'h00, 8'ha0, 8'he0, 8'h00, 8'h00, 8'hc0, 8'h00, 8'h00, 8'h00, 8'hc0,
    8'h20, 8'h00, 8'h00, 8'hc0, 8'h40, 8'h00, 8'h00, 8'hc0, 8'h60, 8'h00, 8'h00, 8'hc0,
    8'h80, 8'h00, 8'h00, 8'hc0, 8'ha0, 8'h00, 8'h00, 8'hc0, 8'hc0, 8'h00, 8'h00, 8'hc0,
    8'he0, 8'h00, 8'h00, 8'he0, 8'h00, 8'h00, 8'h00, 8'he0, 8'h20, 8'h00, 8'h00, 8'he0,
    8'h40, 8'h00, 8'h00, 8'he0, 8'h60, 8'h00, 8'h00, 8'he0, 8'h80, 8'h00, 8'h00, 8'he0,
    8'ha0, 8'h00, 8'h00, 8'he0, 8'hc0, 8'h00, 8'h00, 8'he0, 8'he0, 8'h00, 8'h40, 8'h00,
    8'h00, 8'h00, 8'h40, 8'h00, 8'h20, 8'h00, 8'h40, 8'h00, 8'h40, 8'h00, 8'h40, 8'h00,
    8'h60, 8'h00, 8'h40, 8'h00, 8'h80, 8'h00, 8'h40, 8'h00, 8'ha0, 8'h00, 8'h40, 8'h00,
    8'hc0, 8'h00, 8'h40, 8'h00, 8'he0, 8'h00, 8'h40, 8'h20, 8'h00, 8'h00, 8'h40, 8'h20,
    8'h20, 8'h00, 8'h40, 8'h20, 8'h40, 8'h00, 8'h40, 8'h20, 8'h60, 8'h00, 8'h40, 8'h20,
    8'h80, 8'h00, 8'h40, 8'h20, 8'ha0, 8'h00, 8'h40, 8'h20, 8'hc0, 8'h00, 8'h40, 8'h20,
    8'he0, 8'h00, 8'h40, 8'h40, 8'h00, 8'h00, 8'h40, 8'h40, 8'h20, 8'h00, 8'h40, 8'h40,
    8'h40, 8'h00, 8'h40, 8'h40, 8'h60, 8'h00, 8'h40, 8'h40, 8'h80, 8'h00, 8'h40, 8'h40,
    8'ha0, 8'h00, 8'h40, 8'h40, 8'hc0, 8'h00, 8'h40, 8'h40, 8'he0, 8'h00, 8'h40, 8'h60,
    8'h00, 8'h00, 8'h40, 8'h60, 8'h20, 8'h00, 8'h40, 8'h60, 8'h40, 8'h00, 8'h40, 8'h60,
    8'h60, 8'h00, 8'h40, 8'h60, 8'h80, 8'h00, 8'h40, 8'h60, 8'ha0, 8'h00, 8'h40, 8'h60,
    8'hc0, 8'h00, 8'h40, 8'h60, 8'he0, 8'h00, 8'h40, 8'h80, 8'h00, 8'h00, 8'h40, 8'h80,
    8'h20, 8'h00, 8'h40, 8'h80, 8'h40, 8'h00, 8'h40, 8'h80, 8'h60, 8'h00, 8'h40, 8'h80,
    8'h80, 8'h00, 8'h40, 8'h80, 8'ha0, 8'h00, 8'h40, 8'h80, 8'hc0, 8'h00, 8'h40, 8'h80,
    8'he0, 8'h00, 8'h40, 8'ha0, 8'h00, 8'h00, 8'h40, 8'ha0, 8'h20, 8'h00, 8'h40, 8'ha0,
    8'h40, 8'h00, 8'h40, 8'ha0, 8'h60, 8'h00, 8'h40, 8'ha0, 8'h80, 8'h00, 8'h40, 8'ha0,
    8'ha0, 8'h00, 8'h40, 8'ha0, 8'hc0, 8'h00, 8'h40, 8'ha0, 8'he0, 8'h00, 8'h40, 8'hc0,
    8'h00, 8'h00, 8'h40, 8'hc0, 8'h20, 8'h00, 8'h40, 8'hc0, 8'h40, 8'h00, 8'h40, 8'hc0,
    8'h60, 8'h00, 8'h40, 8'hc0, 8'h80, 8'h00, 8'h40, 8'hc0, 8'ha0, 8'h00, 8'h40, 8'hc0,
    8'hc0, 8'h00, 8'h40, 8'hc0, 8'he0, 8'h00, 8'h40, 8'he0, 8'h00, 8'h00, 8'h40, 8'he0,
    8'h20, 8'h00, 8'h40, 8'he0, 8'h40, 8'h00, 8'h40, 8'he0, 8'h60, 8'h00, 8'h40, 8'he0,
    8'h80, 8'h00, 8'h40, 8'he0, 8'ha0, 8'h00, 8'h40, 8'he0, 8'hc0, 8'h00, 8'h40, 8'he0,
    8'he0, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h80, 8'h00, 8'h20, 8'h00, 8'h80, 8'h00,
    8'h40, 8'h00, 8'h80, 8'h00, 8'h60, 8'h00, 8'h80, 8'h00, 8'h80, 8'h00, 8'h80, 8'h00,
    8'ha0, 8'h00, 8'h80, 8'h00, 8'hc0, 8'h00, 8'h80, 8'h00, 8'he0, 8'h00, 8'h80, 8'h20,
    8'h00, 8'h00, 8'h80, 8'h20, 8'h20, 8'h00, 8'h80, 8'h20, 8'h40, 8'h00, 8'h80, 8'h20,
    8'h60, 8'h00, 8'h80, 8'h20, 8'h80, 8'h00, 8'h80, 8'h20, 8'ha0, 8'h00, 8'h80, 8'h20,
    8'hc0, 8'h00, 8'h80, 8'h20, 8'he0, 8'h00, 8'h80, 8'h40, 8'h00, 8'h00, 8'h80, 8'h40,
    8'h20, 8'h00, 8'h80, 8'h40, 8'h40, 8'h00, 8'h80, 8'h40, 8'h60, 8'h00, 8'h80, 8'h40,
    8'h80, 8'h00, 8'h80, 8'h40, 8'ha0, 8'h00, 8'h80, 8'h40, 8'hc0, 8'h00, 8'h80, 8'h40,
    8'he0, 8'h00, 8'h80, 8'h60, 8'h00, 8'h00, 8'h80, 8'h60, 8'h20, 8'h00, 8'h80, 8'h60,
    8'h40, 8'h00, 8'h80, 8'h60, 8'h60, 8'h00, 8'h80, 8'h60, 8'h80, 8'h00, 8'h80, 8'h60,
    8'ha0, 8'h00, 8'h80, 8'h60, 8'hc0, 8'h00, 8'h80, 8'h60, 8'he0, 8'h00, 8'h80, 8'h80,
    8'h00, 8'h00, 8'h80, 8'h80, 8'h20, 8'h00, 8'h80, 8'h80, 8'h40, 8'h00, 8'h80, 8'h80,
    8'h60, 8'h00, 8'h80, 8'h80, 8'h80, 8'h00, 8'h80, 8'h80, 8'ha0, 8'h00, 8'h80, 8'h80,
    8'hc0, 8'h00, 8'h80, 8'h80, 8'he0, 8'h00, 8'h80, 8'ha0, 8'h00, 8'h00, 8'h80, 8'ha0,
    8'h20, 8'h00, 8'h80, 8'ha0, 8'h40, 8'h00, 8'h80, 8'ha0, 8'h60, 8'h00, 8'h80, 8'ha0,
    8'h80, 8'h00, 8'h80, 8'ha0, 8'ha0, 8'h00, 8'h80, 8'ha0, 8'hc0, 8'h00, 8'h80, 8'ha0,
    8'he0, 8'h00, 8'h80, 8'hc0, 8'h00, 8'h00, 8'h80, 8'hc0, 8'h20, 8'h00, 8'h80, 8'hc0,
    8'h40, 8'h00, 8'h80, 8'hc0, 8'h60, 8'h00, 8'h80, 8'hc0, 8'h80, 8'h00, 8'h80, 8'hc0,
    8'ha0, 8'h00, 8'h80, 8'hc0, 8'hc0, 8'h00, 8'h80, 8'hc0, 8'he0, 8'h00, 8'h80, 8'he0,
    8'h00, 8'h00, 8'h80, 8'he0, 8'h20, 8'h00, 8'h80, 8'he0, 8'h40, 8'h00, 8'h80, 8'he0,
    8'h60, 8'h00, 8'h80, 8'he0, 8'h80, 8'h00, 8'h80, 8'he0, 8'ha0, 8'h00, 8'h80, 8'he0,
    8'hc0, 8'h00, 8'h80, 8'he0, 8'he0, 8'h00, 8'hc0, 8'h00, 8'h00, 8'h00, 8'hc0, 8'h00,
    8'h20, 8'h00, 8'hc0, 8'h00, 8'h40, 8'h00, 8'hc0, 8'h00, 8'h60, 8'h00, 8'hc0, 8'h00,
    8'h80, 8'h00, 8'hc0, 8'h00, 8'ha0, 8'h00, 8'hc0, 8'h00, 8'hc0, 8'h00, 8'hc0, 8'h00,
    8'he0, 8'h00, 8'hc0, 8'h20, 8'h00, 8'h00, 8'hc0, 8'h20, 8'h20, 8'h00, 8'hc0, 8'h20,
    8'h40, 8'h00, 8'hc0, 8'h20, 8'h60, 8'h00, 8'hc0, 8'h20, 8'h80, 8'h00, 8'hc0, 8'h20,
    8'ha0, 8'h00, 8'hc0, 8'h20, 8'hc0, 8'h00, 8'hc0, 8'h20, 8'he0, 8'h00, 8'hc0, 8'h40,
    8'h00, 8'h00, 8'hc0, 8'h40, 8'h20, 8'h00, 8'hc0, 8'h40, 8'h40, 8'h00, 8'hc0, 8'h40,
    8'h60, 8'h00, 8'hc0, 8'h40, 8'h80, 8'h00, 8'hc0, 8'h40, 8'ha0, 8'h00, 8'hc0, 8'h40,
    8'hc0, 8'h00, 8'hc0, 8'h40, 8'he0, 8'h00, 8'hc0, 8'h60, 8'h00, 8'h00, 8'hc0, 8'h60,
    8'h20, 8'h00, 8'hc0, 8'h60, 8'h40, 8'h00, 8'hc0, 8'h60, 8'h60, 8'h00, 8'hc0, 8'h60,
    8'h80, 8'h00, 8'hc0, 8'h60, 8'ha0, 8'h00, 8'hc0, 8'h60, 8'hc0, 8'h00, 8'hc0, 8'h60,
    8'he0, 8'h00, 8'hc0, 8'h80, 8'h00, 8'h00, 8'hc0, 8'h80, 8'h20, 8'h00, 8'hc0, 8'h80,
    8'h40, 8'h00, 8'hc0, 8'h80, 8'h60, 8'h00, 8'hc0, 8'h80, 8'h80, 8'h00, 8'hc0, 8'h80,
    8'ha0, 8'h00, 8'hc0, 8'h80, 8'hc0, 8'h00, 8'hc0, 8'h80, 8'he0, 8'h00, 8'hc0, 8'ha0,
    8'h00, 8'h00, 8'hc0, 8'ha0, 8'h20, 8'h00, 8'hc0, 8'ha0, 8'h40, 8'h00, 8'hc0, 8'ha0,
    8'h60, 8'h00, 8'hc0, 8'ha0, 8'h80, 8'h00, 8'hc0, 8'ha0, 8'ha0, 8'h00, 8'hc0, 8'ha0,
    8'hc0, 8'h00, 8'hc0, 8'ha0, 8'he0, 8'h00, 8'hc0, 8'hc0, 8'h00, 8'h00, 8'hc0, 8'hc0,
    8'h20, 8'h00, 8'hc0, 8'hc0, 8'h40, 8'h00, 8'hc0, 8'hc0, 8'h60, 8'h00, 8'hc0, 8'hc0,
    8'h80, 8'h00, 8'hc0, 8'hc0, 8'ha0, 8'h00, 8'hf0, 8'hfb, 8'hff, 8'h00, 8'ha4, 8'ha0,
    8'ha0, 8'h00, 8'h80, 8'h80, 8'h80, 8'h00, 8'h00, 8'h00, 8'hff, 8'h00, 8'h00, 8'hff,
    8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'h00, 8'hff, 8'h00, 8'h00, 8'h00, 8'hff, 8'h00,
    8'hff, 8'h00, 8'hff, 8'hff, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'h00
};

`endif